/* encoding :utf-8  实例数组*/
module top_module(
           input [399:0] a, b,
           input cin,
           output cout,
           output [399:0] sum );

wire [99:0] intermediate_cin,intermediate_cout;

bcd_fadd u_bcd_fadd[99:0](
             a[399:0],
             b[399:0],
             intermediate_cin[99:0],
             intermediate_cout[99:0],
             sum[399:0]
         );

assign intermediate_cin[0] = cin;
assign intermediate_cin[99:1] = intermediate_cout[98:0];
assign cout = intermediate_cout[99];
endmodule

    /*
    module top_module(
            input [399:0] a, b,
            input cin,
            output cout,
            output [399:0] sum );
     
    wire [99:0] cout_temp;
     
    bcd_fadd u_bcd_fadd(
                 .a(a[3:0]),
                 .b(b[3:0]),
                 .cin(cin),
                 .cout(cout_temp[0]),
                 .sum(sum[3:0])
             );
    generate
        genvar i;
        for(i=1; i<100; i=i+1) begin : block1
            bcd_fadd u_bcd_fadd(
                         .a(a[4*i+3 : 4*i]),
                         .b(b[4*i+3 : 4*i]),
                         .cin(cout_temp[i-1]),
                         .cout(cout_temp[i]),
                         .sum(sum[4*i+3 : 4*i])
                     );
        end
    endgenerate
    assign cout = cout_temp[99];
    endmodule
    */
